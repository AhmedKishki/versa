    // Each of the 14 bits in the binary pattern corresponds to a specific segment.
    // Each segment can be turned ON or OFF by setting its corresponding bit in the 14-bit pattern.
    localparam pat_len = 52;
    wire [13:0] display_pat[0:pat_len-1];
    assign display_pat[0] = 14'b10001000110110;  // H
    assign display_pat[1] = 14'b10000000111001;  // E
    assign display_pat[2] = 14'b00000000111000;  // L
    assign display_pat[3] = 14'b00000000111000;  // L
    assign display_pat[4] = 14'b00000000111111;  // O
    assign display_pat[5] = 14'b00000000000000;
    assign display_pat[6] = 14'b01010000110110;  // W
    assign display_pat[7] = 14'b00000000111111;  // O
    assign display_pat[8] = 14'b10010100110001;  // R
    assign display_pat[9] = 14'b00000000111000;  // L
    assign display_pat[10] = 14'b01000001110000;  // D
    assign display_pat[11] = 14'b00000000000000;
    assign display_pat[12] = 14'b10000000110001;  // F
    assign display_pat[13] = 14'b10010100110001;  // R
    assign display_pat[14] = 14'b00000000111111;  // O
    assign display_pat[15] = 14'b00000101110110;  // M
    assign display_pat[16] = 14'b00000000000000;
    assign display_pat[17] = 14'b10001000110011;  // P
    assign display_pat[18] = 14'b10010100110001;  // R
    assign display_pat[19] = 14'b00000000111111;  // O
    assign display_pat[20] = 14'b00000000001110;  // J
    assign display_pat[21] = 14'b10000000111001;  // E
    assign display_pat[22] = 14'b00000000111001;  // C
    assign display_pat[23] = 14'b00100010000001;  // T
    assign display_pat[24] = 14'b00000000000000;
    assign display_pat[25] = 14'b00100010000001;  // T
    assign display_pat[26] = 14'b10010100110001;  // R
    assign display_pat[27] = 14'b10000000111001;  // E
    assign display_pat[28] = 14'b00000000111000;  // L
    assign display_pat[29] = 14'b00000000111000;  // L
    assign display_pat[30] = 14'b00100010001001;  // I
    assign display_pat[31] = 14'b10001000101101;  // S
    assign display_pat[32] = 14'b00000000000000;
    assign display_pat[33] = 14'b00000000111111;  // O
    assign display_pat[34] = 14'b00010001110110;  // N
    assign display_pat[35] = 14'b00000000000000;
    assign display_pat[36] = 14'b00100010000001;  // T
    assign display_pat[37] = 14'b10001000110110;  // H
    assign display_pat[38] = 14'b10000000111001;  // E
    assign display_pat[39] = 14'b00000000000000;
    assign display_pat[40] = 14'b01000100110000;  // V
    assign display_pat[41] = 14'b10000000111001;  // E
    assign display_pat[42] = 14'b10010100110001;  // R
    assign display_pat[43] = 14'b10001000101101;  // S
    assign display_pat[44] = 14'b10001000110111;  // A
    assign display_pat[45] = 14'b00000000000000;
    assign display_pat[46] = 14'b10010100111001;  // B
    assign display_pat[47] = 14'b00000000111111;  // O
    assign display_pat[48] = 14'b10001000110111;  // A
    assign display_pat[49] = 14'b10010100110001;  // R
    assign display_pat[50] = 14'b01000001110000;  // D
    assign display_pat[51] = 14'b00000000000000;
